----------------------------------------------------------------------
--! @file  
--! @brief 
--!
--!
--! @author 
--! @date 
--! @version  
--! 
-- note 
--! @todo 
--! @test 
--! @bug  
--!
----------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pulse_integrator is
	port (
		isl_clk50Mhz : in std_logic;
		rst : in std_logic
	);
end entity pulse_integrator;

architecture RTL of pulse_integrator is
	
begin

end architecture RTL;
