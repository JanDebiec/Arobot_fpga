--! @mainpage notitle
--!
--! additional information about arobot fpga copy from msystem, TO BE EDITED
--!
--! @TODO: change the content of arobot doxy
--! @tableofcontents
--! @section  structure
--! @subsection  H2F_interface
--!
--! | interface    | functionality   | top-file name            |
--! |:------------:|:---------------:|:------------------------:|
--! | light-weight | @ref h2flw_addr | arobot_constant_pkg.vhd |
--!
--!
--!
--! @section  formal
--!
--! | item    | functionality   | top-file name            |
--! |:------------:|:---------------:|:------------------------:|
--! | version | @ref fpga_version | version.vhd |
--! | style guide | @ref style_guide | doxy_styleguide.vhd |



